class axi4lite_test extends uvm_test;

  `uvm_component_utils(axi4lite_test)
  
  axi4lite_env  env;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction 

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    env = axi4lite_env::type_id::create("env",this);
  endfunction

  virtual task run_phase(uvm_phase phase); 
 
    axi4lite_sequence seq; 

  
    super.run_phase(phase);
    
    phase.raise_objection(this);

    seq = axi4lite_sequence::type_id::create("seq");
    seq.start(env.agent.sequencer);
    
    phase.drop_objection(this);
  endtask 

endclass